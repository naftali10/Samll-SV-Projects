`include "defines.sv"
