`include "defines.sv"
`include "naive_FSM.sv"
