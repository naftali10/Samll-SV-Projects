`define WINDOW_SZ 128
`define PATTERN_SZ 8
`define PATTERN `PATTERN_SZ'he8
`define SR_SZ 8
`define OUT_SZ 8
